`define _CACHE_SIZE 'd1
`define _CACHE_TYPE x

`define _CACHE_TYPE_DATA 'd0
`define _DATA_CACHE_SIZE 'h100
`define _DATA_CACHE_PAYLOAD mem_cell[0] <= 1; \
                            mem_cell[0] <= 1; \
                            mem_cell[0] <= 1;
`define _CACHE_TYPE_INST 'd1
`define _INST_CACHE_SIZE 'h1ec
`define _INST_CACHE_PAYLOAD mem_cell[0] <= 1; \
                            mem_cell[0] <= 1; \
                            mem_cell[0] <= 1;



