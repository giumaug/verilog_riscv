`define _CACHE_SIZE 1
`define _CACHE_PAYLOAD_SIZE 1
`define _CACHE_PAYLOAD {8'd0, 8'd1,8'd0, 8'd1,8'd0, 8'd1,8'd0, 8'd1}
`define __CACHE_PAYLOAD 1

`define _DATA_CACHE_SIZE 0x100
`define _DATA_CACHE_PAYLOAD_SIZE 0x1c
`define _DATA_CACHE_PAYLOAD {16'd4, 16'd4}

`define _INST_CACHE_SIZE
`define _INST_CACHE_PAYLOAD_SIZE
`define _INST_CACHE_PAYLOAD



