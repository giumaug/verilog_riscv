`define CACHE_SIZE 0x1
`define CACHE_PAYLOAD_SIZE 0x1
`define CACHE_PAYLOAD {8'd0}

`define DATA_CACHE_SIZE 0x100
`define DATA_CACHE_PAYLOAD_SIZE 0x1c
`define DATA_CACHE_PAYLOAD {16'd4, 16'd4}

`define INST_CACHE_SIZE
`define INST_CACHE_PAYLOAD_SIZE
`define INST_CACHE_PAYLOAD



