module memory_controller(input[31:0] address_1,
                         input[31:0] i_val_1,
                         input op_type_1,
					     input[31:0] address_2,
                         input[31:0] i_val_2,
                         input op_type_2,
                         output[31:0] o_val_1,
						 output[31:0] o_val_2);

	always @(...)
    begin

	end
endmodule     
